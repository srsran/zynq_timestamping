library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library UNISIM;
use UNISIM.vcomponents.all;

entity single_port_memory is
  generic (
    g_MEM_CLOCK_DOMAIN_TYPE: string := "INDEPENDENT"; --! Read/write clock domain type. Supported types: "INDEPENDENT".
    g_MEM_TYPE : string := "ramb36e2"; --! Memory instantiation type. Supported types: "**ramb36e2**", "**ramb36e1**"
    g_DATA_WIDTH : integer := 32; --! Memory data bus width.
    g_ADDRESS_WIDTH : integer := 15 --! Memory size E.g. g_ADDRESS_WIDTH=15 -> 2^15 words.
  );
  port (
    rd_clk   : in std_logic; --! Read clock.
    wr_clk   : in std_logic; --! Write clock.

    rd_reset : in std_logic; --! Active hight read reset (@rd_clk).
    wr_reset : in std_logic; --! Active hight write reset (@wr_clk).

    wr_address : in std_logic_vector(g_ADDRESS_WIDTH-1 downto 0); --! Write address (@wr_clk).
    wr_din : in std_logic_vector(g_DATA_WIDTH-1 downto 0); --! Write data in (@wr_clk).
    wr_byte_wide : in std_logic_vector(7 downto 0); --! Write byte wide (@wr_clk).
    wr_enable : in std_logic; --! Write enable (@wr_clk).

    rd_address : in std_logic_vector(g_ADDRESS_WIDTH-1 downto 0); --! Read address (@rd_clk) .
    rd_dout : out std_logic_vector(g_DATA_WIDTH-1 downto 0); --! Read data out (@rd_clk).
    rd_enable : in std_logic --! Read enable (@rd_clk).
  );
end entity;

architecture rtl of single_port_memory is

  -- **********************************
  -- definition of constants
  -- **********************************

  -- RAMB instantiation constants
  constant cnt_RAMB_parity_width : integer := integer(g_DATA_WIDTH / 8);  -- 1 parity bit per byte
  constant cnt_RAMB_data_width : integer := g_DATA_WIDTH + cnt_RAMB_parity_width;

  -- **********************************
  -- internal signals
  -- **********************************

  -- RAMB instantiation signals
  signal wr_address_s : std_logic_vector(15 downto 0):=(others => '0');
  signal wr_din_s : std_logic_vector(31 downto 0):=(others => '0');
  signal rd_address_s : std_logic_vector(15 downto 0):=(others => '0');
  signal rd_dout_s : std_logic_vector(31 downto 0):=(others => '0');

begin

  -- map signals and ports
  wr_address_s(g_ADDRESS_WIDTH-1 downto 0) <= wr_address;
  wr_din_s(g_DATA_WIDTH-1 downto 0) <= wr_din;
  rd_address_s(g_ADDRESS_WIDTH-1 downto 0) <= rd_address;
  rd_dout <= rd_dout_s(g_DATA_WIDTH-1 downto 0);

  ramb36e2_gen : if g_MEM_TYPE = "ramb36e2" generate
    ramb36e2_inst : RAMB36E2
      GENERIC MAP (
        -- CASCADE_ORDER_A, CASCADE_ORDER_B: "FIRST", "MIDDLE", "LAST", "NONE"
        CASCADE_ORDER_A => "NONE",
        CASCADE_ORDER_B => "NONE",
        -- CLOCK_DOMAINS: "COMMON", "INDEPENDENT"
        CLOCK_DOMAINS => g_MEM_CLOCK_DOMAIN_TYPE,
        DOB_REG => 1,
        -- Collision check: "ALL", "GENERATE_X_ONLY", "NONE", "WARNING_ONLY"
        SIM_COLLISION_CHECK => "ALL",
        -- DOA_REG, DOB_REG: Optional output register (0, 1)
        DOA_REG => 1,
        -- ENADDRENA/ENADDRENB: Address enable pin enable, "TRUE", "FALSE"
        ENADDRENA => "FALSE",
        ENADDRENB => "FALSE",
        -- EN_ECC_PIPE: ECC pipeline register, "TRUE"/"FALSE"
        EN_ECC_PIPE => "FALSE",
        -- EN_ECC_READ: Enable ECC decoder, "TRUE"/"FALSE"
        EN_ECC_READ => "FALSE",
        -- EN_ECC_WRITE: Enable ECC encoder, "TRUE"/"FALSE"
        EN_ECC_WRITE => "FALSE",
        -- Programmable inversion Attributes: Specifies the use of the built-in programmable inversion
        IS_CLKARDCLK_INVERTED => '0',
        IS_CLKBWRCLK_INVERTED => '0',
        IS_ENARDEN_INVERTED => '0',
        IS_ENBWREN_INVERTED => '0',
        IS_RSTRAMARSTRAM_INVERTED => '0',
        IS_RSTRAMB_INVERTED => '0',
        IS_RSTREGARSTREG_INVERTED => '0',
        IS_RSTREGB_INVERTED => '0',
        -- RDADDRCHANGE: Disable memory access when output value does not change ("TRUE", "FALSE")
        RDADDRCHANGEA => "FALSE",
        RDADDRCHANGEB => "FALSE",
        -- READ_WIDTH_A/B, WRITE_WIDTH_A/B: Read/write width per port
        READ_WIDTH_A => cnt_RAMB_data_width,   -- [0,1,2,4,9,18,36,72]; * since the memory is used as a SDP, then port A is the read port *
        READ_WIDTH_B => 0,                     -- [0,1,2,4,9,18,36,72]
        WRITE_WIDTH_A => 0,                    -- [0,1,2,4,9,18,36,72]
        WRITE_WIDTH_B => cnt_RAMB_data_width,  -- [0,1,2,4,9,18,36,72]; * since the memory is used as a SDP, then port B is the write port *
        -- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG", "REGCE")
        RSTREG_PRIORITY_A => "RSTREG",
        RSTREG_PRIORITY_B => "RSTREG",
        -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_A => X"000000000",
        SRVAL_B => X"000000000",
        -- Sleep Async: Sleep function asynchronous or synchronous ("TRUE", "FALSE")
        SLEEP_ASYNC => "FALSE",
        -- WriteMode: "WRITE_FIRST", "NO_CHANGE", "READ_FIRST"
        WRITE_MODE_A => "NO_CHANGE",
        WRITE_MODE_B => "NO_CHANGE",
        -- INIT_A, INIT_B: Initial values on output ports
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        -- Initialization File: RAM initialization file
        INIT_FILE => "NONE",
        -- INIT_00 to INIT_7F: Initial contents of data memory array
        INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
        -- INITP_00 to INITP_0F: Initial contents of parity memory array
        INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
      )
    PORT MAP (
      -- Cascade Signals outputs: Multi-BRAM cascade signals
      CASDOUTA => OPEN,                                       -- ** NOT USED ** 32-bit output: Port A cascade output data
      CASDOUTB => OPEN,                                       -- ** NOT USED ** 32-bit output: Port B cascade output data
      CASDOUTPA => OPEN,                                      -- ** NOT USED ** 4-bit output: Port A cascade output parity data
      CASDOUTPB => OPEN,                                      -- ** NOT USED ** 4-bit output: Port B cascade output parity data
      CASOUTDBITERR => OPEN,                                  -- ** NOT USED ** 1-bit output: DBITERR cascade output
      CASOUTSBITERR => OPEN,                                  -- ** NOT USED ** 1-bit output: SBITERR cascade output
      -- ECC Signals outputs: Error Correction Circuitry ports
      DBITERR => OPEN,                                        -- ** NOT USED ** 1-bit output: Double bit error status
      ECCPARITY => OPEN,                                      -- ** NOT USED ** 8-bit output: Generated error correction parity
      RDADDRECC => OPEN,                                      -- ** NOT USED ** 9-bit output: ECC Read Address
      SBITERR => OPEN,                                        -- ** NOT USED ** 1-bit output: Single bit error status
      -- Port A Data outputs: Port A data
      DOUTADOUT => rd_dout_s,                                 -- 32-bit output: Port A data/LSB data; * since the memory is used as a SDP, then port A is the read port *
      DOUTPADOUTP => OPEN,                                    -- ** NOT USED ** 4-bit output: Port A parity/LSB parity
      -- Port B Data outputs: Port B data
      DOUTBDOUT => OPEN,                                      -- ** NOT USED ** 32-bit output: Port B data/MSB data; * since the memory is used as a SDP, then port B is the write port *
      DOUTPBDOUTP => OPEN,                                    -- ** NOT USED ** @TO_BE_TESTED: this extra 4 bits might be useful in the future; 4-bit output: Port B parity/MSB parity
      -- Cascade Signals inputs: Multi-BRAM cascade signals
      CASDIMUXA => '0',                                       -- ** NOT USED (initialized accordging to table 1-12 [UG573])** 1-bit input: Port A input data (0=DINA, 1=CASDINA)
      CASDIMUXB => '0',                                       -- ** NOT USED (initialized accordging to table 1-12 [UG573])** 1-bit input: Port B input data (0=DINB, 1=CASDINB)
      CASDINA => (others => '0'),                             -- ** NOT USED ** 32-bit input: Port A cascade input data
      CASDINB => (others => '0'),                             -- ** NOT USED ** 32-bit input: Port B cascade input data
      CASDINPA => (others => '0'),                            -- ** NOT USED ** 4-bit input: Port A cascade input parity data
      CASDINPB => (others => '0'),                            -- ** NOT USED ** 4-bit input: Port B cascade input parity data
      CASDOMUXA => '0',                                       -- ** NOT USED (initialized accordging to table 1-12 [UG573])** 1-bit input: Port A unregistered data (0=BRAM data, 1=CASDINA)
      CASDOMUXB => '0',                                       -- ** NOT USED (initialized accordging to table 1-12 [UG573])** 1-bit input: Port B unregistered data (0=BRAM data, 1=CASDINB)
      CASDOMUXEN_A => '1',                                    -- ** NOT USED (initialized accordging to table 1-12 [UG573])** 1-bit input: Port A unregistered output data enable
      CASDOMUXEN_B => '1',                                    -- ** NOT USED (initialized accordging to table 1-12 [UG573])** 1-bit input: Port B unregistered output data enable
      CASINDBITERR => '0',                                    -- ** NOT USED ** 1-bit input: DBITERR cascade input
      CASINSBITERR => '0',                                    -- ** NOT USED ** 1-bit input: SBITERR cascade input
      CASOREGIMUXA => '0',                                    -- ** NOT USED (initialized accordging to table 1-12 [UG573])** 1-bit input: Port A registered data (0=BRAM data, 1=CASDINA)
      CASOREGIMUXB => '0',                                    -- ** NOT USED (initialized accordging to table 1-12 [UG573])** 1-bit input: Port B registered data (0=BRAM data, 1=CASDINB)
      CASOREGIMUXEN_A => '1',                                 -- ** NOT USED (initialized accordging to table 1-12 [UG573])** 1-bit input: Port A registered output data enable
      CASOREGIMUXEN_B => '1',                                 -- ** NOT USED (initialized accordging to table 1-12 [UG573])** 1-bit input: Port B registered output data enable
      -- ECC Signals inputs: Error Correction Circuitry ports
      ECCPIPECE => '0',                                       -- ** NOT USED ** 1-bit input: ECC Pipeline Register Enable
      INJECTDBITERR => '0',                                   -- ** NOT USED (initialized accordging to table 1-12 [UG573])** 1-bit input: inject a double bit error
      INJECTSBITERR => '0',                                   -- ** NOT USED (initialized accordging to table 1-12 [UG573])** 1-bit input: inject a single bit error
      -- Port A Address/Control Signals inputs: Port A address and control signals
      ADDRARDADDR => rd_address_s(14 downto 0),               -- 15-bit input: A/Read port address; * since the memory is used as a SDP, then port A is the read port *
      ADDRENA => '1',                                         -- 1-bit input: Active-High A/Read port address enable
      CLKARDCLK => rd_clk,                                    -- 1-bit input: A/Read port clock
      ENARDEN => rd_enable,                                   -- 1-bit input: Port A enable/Read enable; * since the memory is used as a SDP, then port A is the read port *
      REGCEAREGCE => '1',                                     -- 1-bit input: Port A register enable/Register enable
      RSTRAMARSTRAM => rd_reset,                              -- 1-bit input: Port A set/reset
      RSTREGARSTREG => rd_reset,                              -- 1-bit input: Port A register set/reset
      SLEEP => '0',                                           -- @TO_BE_TESTED: in the future it might be interesting to be able to power-off part of the logic; 1-bit input: Sleep Mode
      WEA => (others => '0'),                                 -- ** NOT USED ** 4-bit input: Port A write enable; * since the memory is used as a SDP, then port A is the read port (and this port is thus not used) *
      -- Port A Data inputs: Port A data
      DINADIN => (others => '0'),                             -- ** NOT USED ** 32-bit input: Port A data/LSB data; * since the memory is used as a SDP, then port A is the read port *
      DINPADINP => (others => '0'),                           -- ** NOT USED ** @TO_BE_TESTED: this extra 4 bits might be useful in the future; 4-bit input: Port A parity/LSB parity
      -- Port B Address/Control Signals inputs: Port B address and control signals
      ADDRBWRADDR => wr_address_s(14 downto 0),               -- 15-bit input: B/Write port address; * since the memory is used as a SDP, then port B is the write port *
      ADDRENB => '1',                                         -- 1-bit input: Active-High B/Write port address enable
      CLKBWRCLK => wr_clk,                                    -- 1-bit input: B/Write port clock
      ENBWREN => wr_enable,                                   -- 1-bit input: Port B enable/Write enable; * since the memory is used as a SDP, then port B is the write port *
      REGCEB => '1',                                          -- 1-bit input: Port B register enable
      RSTRAMB => wr_reset,                                    -- 1-bit input: Port B set/reset
      RSTREGB => wr_reset,                                    -- 1-bit input: Port B register set/reset
      WEBWE => wr_byte_wide,                                  -- 8-bit input: Port B write enable/Write enable; * since the memory is used as a SDP, then port B is the write port *
      -- Port B Data inputs: Port B data
      DINBDIN => wr_din_s,                                    -- 32-bit input: Port B data/MSB data; * since the memory is used as a SDP, then port B is the write port *
      DINPBDINP => (others => '0')                            -- ** NOUT USED ** 4-bit input: Port B parity/MSB parity
    );
  end generate ramb36e2_gen;

  ramb36e1_gen : if g_MEM_TYPE = "ramb36e1" generate
    ramb36e1_inst : RAMB36E1
      GENERIC MAP (
        -- Collision check: "ALL", "GENERATE_X_ONLY", "NONE", "WARNING_ONLY"
        SIM_COLLISION_CHECK => "ALL",
        -- DOA_REG, DOB_REG: Optional output register (0, 1)
        DOA_REG => 1,
        DOB_REG => 1,
        -- Error Correction Circuitry (ECC): Encoder/decoder enable (TRUE/FALSE)
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_A => "NONE",
        RAM_EXTENSION_B => "NONE",
        RAM_MODE => "TDP", -- "SDP" (Single Dual Port) or "TDP" (True Dual Port)
        --RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE", -- "PERFORMANCE" or "DELAYED_WRITE"
        -- READ_WIDTH_A/B, WRITE_WIDTH_A/B: Read/write width per port
        READ_WIDTH_A => cnt_RAMB_data_width,   -- [0,1,2,4,9,18,36,72]; * since the memory is used as a SDP, then port A is the read port *
        READ_WIDTH_B => 0,                     -- [0,1,2,4,9,18,36,72]
        WRITE_WIDTH_A => 0,                    -- [0,1,2,4,9,18,36,72]
        WRITE_WIDTH_B => cnt_RAMB_data_width,  -- [0,1,2,4,9,18,36,72]; * since the memory is used as a SDP, then port B is the write port *
        -- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG", "REGCE")
        RSTREG_PRIORITY_A => "RSTREG",
        RSTREG_PRIORITY_B => "RSTREG",
        -- WriteMode: "WRITE_FIRST", "NO_CHANGE", "READ_FIRST"
        WRITE_MODE_A => "WRITE_FIRST",  -- according to UG473 p.21, only WF and RF are supported in SDP mode
        WRITE_MODE_B => "WRITE_FIRST",  -- according to UG473 p.21, only WF and RF are supported in SDP mode
        -- Simulation Device: Must be set to "7SERIES" for simulation behavior
        SIM_DEVICE => "7SERIES",
        INIT_FILE => "NONE",
        -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_A => X"000000000",
        SRVAL_B => X"000000000",
        -- INIT_A, INIT_B: Initial values on output ports
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        -- INIT_00 to INIT_7F: Initial contents of data memory array
        INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
        -- INITP_00 to INITP_0F: Initial contents of parity memory array
        INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
      )
    PORT MAP (
      -- Cascade Signals outputs: Multi-BRAM cascade signals
      CASCADEOUTA => OPEN,                                    -- ** NOT USED ** 1-bit A port cascade output
      CASCADEOUTB => OPEN,                                    -- ** NOT USED ** 1-bit B port cascade output
      -- ECC Signals: 1-bit (each) Error Correction Circuitry ports
      DBITERR => OPEN,                                        -- ** NOT USED ** 1-bit double bit error status output
      ECCPARITY => OPEN,                                      -- ** NOT USED ** 8-bit generated error correction parity
      RDADDRECC => OPEN,                                      -- ** NOT USED ** 9-bit ECC read address
      SBITERR => OPEN,                                        -- ** NOT USED ** 1-bit Single bit error status output
      -- Port A Data outputs: Port A data
      DOADO => rd_dout_s,                                     -- 32-bit output: Port A data/LSB data; * since the memory is used as a SDP, then port A is the read port *
      DOPADOP => OPEN,                                        -- ** NOT USED ** 4-bit output: Port A parity/LSB parity; * the parity bits are used to carry the DAC valid and enable signals *
      -- Port B Data outputs: Port B data
      DOBDO => OPEN,                                          -- ** NOT USED ** 32-bit output: Port B data/MSB data; * since the memory is used as a SDP, then port B is the write port *
      DOPBDOP => OPEN,                                        -- ** NOT USED ** @TO_BE_TESTED: this extra 4 bits might be useful in the future; 4-bit output: Port B parity/MSB parity
      -- Cascade Signals inputs: Multi-BRAM cascade signals
      -- Cascade Signals: 1-bit (each) BRAM cascade ports (to create 72kx1)
      CASCADEINA => '0',                                      -- 1-bit A port cascade input
      CASCADEINB => '0',                                      -- 1-bit B port cascade input
      -- ECC Signals: 1-bit (each) Error Correction Circuitry ports
      INJECTDBITERR => '0',                                   -- 1-bit Inject a double bit error
      INJECTSBITERR => '0',                                   -- 1-bit Inject a single bit error                                   -- ** NOT USED (initialized accordging to table 1-12 [UG573])** 1-bit input: inject a single bit error
      -- Port A Address/Control Signals inputs: Port A address and control signals
      ADDRARDADDR => rd_address_s,                            -- 16-bit input: A/Read port address; * since the memory is used as a SDP, then port A is the read port *
      CLKARDCLK => rd_clk,                                    -- 1-bit input: A/Read port clock
      ENARDEN => rd_enable,                                   -- 1-bit input: Port A enable/Read enable; * since the memory is used as a SDP, then port A is the read port *
      REGCEAREGCE => '1',                                     -- 1-bit input: Port A register enable/Register enable
      RSTRAMARSTRAM => rd_reset,                              -- 1-bit input: Port A set/reset
      RSTREGARSTREG => rd_reset,                              -- 1-bit input: Port A register set/reset
      WEA => (others => '0'),                                 -- 4-bit input: Port A write enable; * since the memory is used as a SDP, then port A is the read port (and this port is thus not used) *
      -- Port A Data inputs: Port A data
      DIADI => (others => '0'),                               -- ** NOT USED ** 32-bit input: Port A data/LSB data; * since the memory is used as a SDP, then port A is the read port *
      DIPADIP => (others => '0'),                             -- ** NOT USED ** @TO_BE_TESTED: this extra 4 bits might be useful in the future; 4-bit input: Port A parity/LSB parity
      -- Port B Address/Control Signals inputs: Port B address and control signals
      ADDRBWRADDR => wr_address_s,                            -- 16-bit input: B/Write port address; * since the memory is used as a SDP, then port B is the write port *
      CLKBWRCLK => wr_clk,                                    -- 1-bit input: B/Write port clock
      ENBWREN => wr_enable,                                   -- 1-bit input: Port B enable/Write enable; * since the memory is used as a SDP, then port B is the write port *
      REGCEB => '1',                                          -- 1-bit input: Port B register enable
      RSTRAMB => wr_reset,                                    -- 1-bit input: Port B set/reset
      RSTREGB => wr_reset,                                    -- 1-bit input: Port B register set/reset
      WEBWE => wr_byte_wide,-- 8-bit input: Port B write enable/Write enable; * since the memory is used as a SDP, then port B is the write port *
      -- Port B Data inputs: Port B data
      DIBDI => wr_din_s,                                      -- 32-bit input: Port B data/MSB data; * since the memory is used as a SDP, then port B is the write port *
      DIPBDIP => (others => '0')                              -- 4-bit input: Port B parity/MSB parity; * the parity bits are used to carry the DAC valid and enable signals *
    );
  end generate ramb36e1_gen;


end architecture;